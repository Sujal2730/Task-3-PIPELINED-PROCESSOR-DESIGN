// pipelined_processor.v

// 1. Program Counter
module program_counter (
    input wire clk,
    input wire reset,
    output reg [3:0] pc
);
    always @(posedge clk or posedge reset) begin
        if (reset)
            pc <= 4'b0000;
        else
            pc <= pc + 1;
    end
endmodule

// 2. Instruction Memory
module instruction_memory (
    input wire [3:0] pc,
    output reg [15:0] instruction
);
    reg [15:0] memory [0:15];

    initial begin
        memory[0] = 16'b0000000100100011; // ADD R1, R2, R3
        memory[1] = 16'b0001001000110100; // SUB R2, R3, R4
        memory[2] = 16'b0010001101000000; // LOAD R3, [R4]
        memory[3] = 16'b0000000100100101; // ADD R1, R2, R5
        memory[4] = 16'b0001001100010001; // SUB R3, R1, R1
        memory[5] = 16'b0000000000000000; // NOP or HALT
    end

    always @(*) begin
        if (pc < 6)
            instruction = memory[pc];
        else
            instruction = 16'b0000000000000000; // default NOP for unused PC values
    end
endmodule


// 3. IF/ID Pipeline Register
module if_id_register (
    input wire clk,
    input wire reset,
    input wire [15:0] instruction_in,
    input wire [3:0] pc_in,
    output reg [15:0] instruction_out,
    output reg [3:0] pc_out
);
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            instruction_out <= 0;
            pc_out <= 0;
        end else begin
            instruction_out <= instruction_in;
            pc_out <= pc_in;
        end
    end
endmodule

// 4. Register File
module register_file (
    input wire clk,
    input wire we,
    input wire [3:0] write_addr,
    input wire [7:0] write_data,
    input wire [3:0] read_addr1,
    input wire [3:0] read_addr2,
    output reg [7:0] read_data1,
    output reg [7:0] read_data2
);
    reg [7:0] registers [0:15];

    always @(posedge clk) begin
        if (we) registers[write_addr] <= write_data;
    end

    always @(*) begin
        read_data1 = registers[read_addr1];
        read_data2 = registers[read_addr2];
    end
endmodule

// 5. ID/EX Pipeline Register
module id_ex_register (
    input wire clk,
    input wire reset,
    input wire [3:0] opcode_in, rd_in, rs1_in, rs2_in,
    input wire [7:0] reg_data1_in, reg_data2_in,
    input wire [3:0] pc_in,
    output reg [3:0] opcode_out, rd_out, rs1_out, rs2_out,
    output reg [7:0] reg_data1_out, reg_data2_out,
    output reg [3:0] pc_out
);
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            opcode_out <= 0; rd_out <= 0; rs1_out <= 0; rs2_out <= 0;
            reg_data1_out <= 0; reg_data2_out <= 0; pc_out <= 0;
        end else begin
            opcode_out <= opcode_in; rd_out <= rd_in;
            rs1_out <= rs1_in; rs2_out <= rs2_in;
            reg_data1_out <= reg_data1_in; reg_data2_out <= reg_data2_in;
            pc_out <= pc_in;
        end
    end
endmodule

// 6. ALU
module alu (
    input wire [3:0] opcode,
    input wire [7:0] op1,
    input wire [7:0] op2,
    output reg [7:0] result
);
    always @(*) begin
        case (opcode)
            4'b0000: result = op1 + op2;
            4'b0001: result = op1 - op2;
            4'b0010: result = op1;  // LOAD uses address from Rs1
            default: result = 0;
        endcase
    end
endmodule

// 7. EX/MEM Register
module ex_mem_register (
    input wire clk,
    input wire reset,
    input wire [3:0] opcode_in, rd_in,
    input wire [7:0] alu_result_in, reg_data2_in,
    output reg [3:0] opcode_out, rd_out,
    output reg [7:0] alu_result_out, reg_data2_out
);
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            opcode_out <= 0; rd_out <= 0;
            alu_result_out <= 0; reg_data2_out <= 0;
        end else begin
            opcode_out <= opcode_in; rd_out <= rd_in;
            alu_result_out <= alu_result_in;
            reg_data2_out <= reg_data2_in;
        end
    end
endmodule

// 8. Data Memory
module data_memory (
    input wire clk,
    input wire mem_read,
    input wire [7:0] address,
    output reg [7:0] data_out
);
    reg [7:0] memory [0:255];

    initial begin
        memory[0] = 8'd10;
        memory[1] = 8'd20;
        memory[2] = 8'd30;
        memory[3] = 8'd40;
    end

    always @(*) begin
        if (mem_read)
            data_out = memory[address];
        else
            data_out = 0;
    end
endmodule

// 9. MEM/WB Register
module mem_wb_register (
    input wire clk,
    input wire reset,
    input wire [3:0] opcode_in, rd_in,
    input wire [7:0] alu_result_in, mem_data_in,
    output reg [3:0] opcode_out, rd_out,
    output reg [7:0] write_data_out
);
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            opcode_out <= 0; rd_out <= 0; write_data_out <= 0;
        end else begin
            opcode_out <= opcode_in; rd_out <= rd_in;
            write_data_out <= (opcode_in == 4'b0010) ? mem_data_in : alu_result_in;
        end
    end
endmodule

// Testbench code

module tb_pipelined_processor;

    reg clk;
    reg reset;

    wire [3:0] pc_wire;
    wire [15:0] instr_wire;
    wire [7:0] alu_wire;

    // Instantiate your top module and connect exposed outputs
    top_module uut (
        .clk(clk),
        .reset(reset),
        .pc_out(pc_wire),
        .instr_out(instr_wire),
        .alu_out(alu_wire)
    );

    // Clock generation: 10ns period
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // Reset and simulation control
    initial begin
    reset = 1;
    #20 reset = 0; // release reset
    #500 $finish;
end


	always @(posedge clk) begin
    $display("Time %0t: PC=%h, Instr=%h, ALU=%h", $time, pc_wire, instr_wire, alu_wire);
end

endmodule



